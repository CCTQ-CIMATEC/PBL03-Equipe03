module imm_gen (

);
endmodule